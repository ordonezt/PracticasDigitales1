----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:19:57 07/05/2018 
-- Design Name: 
-- Module Name:    TestMyAnd - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TestMyAnd is
	
	Port	(	a:	in	STD_LOGIC;
				b:	in	STD_LOGIC;
				z:	out STD_LOGIC
			);
			
end TestMyAnd;

architecture Behavioral of TestMyAnd is

begin

	z	<= a AND b;

end Behavioral;

